module ram ( 
	input clk, rst_n,
	input wire [6:0] addr,
	input wire [8:0] data,
	input wire wr_en,
	output reg [8:0] q
);

reg [127:0] reg_sel;
wire [127:0] wr_sel;

reg [8:0] addr_00, addr_01, addr_02, addr_03, addr_04, addr_05, addr_06, addr_07, addr_08, addr_09, addr_0a, addr_0b, addr_0c, addr_0d, addr_0e, addr_0f;
reg [8:0] addr_10, addr_11, addr_12, addr_13, addr_14, addr_15, addr_16, addr_17, addr_18, addr_19, addr_1a, addr_1b, addr_1c, addr_1d, addr_1e, addr_1f;
reg [8:0] addr_20, addr_21, addr_22, addr_23, addr_24, addr_25, addr_26, addr_27, addr_28, addr_29, addr_2a, addr_2b, addr_2c, addr_2d, addr_2e, addr_2f;
reg [8:0] addr_30, addr_31, addr_32, addr_33, addr_34, addr_35, addr_36, addr_37, addr_38, addr_39, addr_3a, addr_3b, addr_3c, addr_3d, addr_3e, addr_3f;
reg [8:0] addr_40, addr_41, addr_42, addr_43, addr_44, addr_45, addr_46, addr_47, addr_48, addr_49, addr_4a, addr_4b, addr_4c, addr_4d, addr_4e, addr_4f;
reg [8:0] addr_50, addr_51, addr_52, addr_53, addr_54, addr_55, addr_56, addr_57, addr_58, addr_59, addr_5a, addr_5b, addr_5c, addr_5d, addr_5e, addr_5f;
reg [8:0] addr_60, addr_61, addr_62, addr_63, addr_64, addr_65, addr_66, addr_67, addr_68, addr_69, addr_6a, addr_6b, addr_6c, addr_6d, addr_6e, addr_6f;
reg [8:0] addr_70, addr_71, addr_72, addr_73, addr_74, addr_75, addr_76, addr_77, addr_78, addr_79, addr_7a, addr_7b, addr_7c, addr_7d, addr_7e, addr_7f;

parameter ADDR_00 = 7'h00;
parameter ADDR_01 = 7'h01;
parameter ADDR_02 = 7'h02;
parameter ADDR_03 = 7'h03;
parameter ADDR_04 = 7'h04;
parameter ADDR_05 = 7'h05;
parameter ADDR_06 = 7'h06;
parameter ADDR_07 = 7'h07;
parameter ADDR_08 = 7'h08;
parameter ADDR_09 = 7'h09;
parameter ADDR_0A = 7'h0A;
parameter ADDR_0B = 7'h0B;
parameter ADDR_0C = 7'h0C;
parameter ADDR_0D = 7'h0D;
parameter ADDR_0E = 7'h0E;
parameter ADDR_0F = 7'h0F;

parameter ADDR_10 = 7'h10;
parameter ADDR_11 = 7'h11;
parameter ADDR_12 = 7'h12;
parameter ADDR_13 = 7'h13;
parameter ADDR_14 = 7'h14;
parameter ADDR_15 = 7'h15;
parameter ADDR_16 = 7'h16;
parameter ADDR_17 = 7'h17;
parameter ADDR_18 = 7'h18;
parameter ADDR_19 = 7'h19;
parameter ADDR_1A = 7'h1A;
parameter ADDR_1B = 7'h1B;
parameter ADDR_1C = 7'h1C;
parameter ADDR_1D = 7'h1D;
parameter ADDR_1E = 7'h1E;
parameter ADDR_1F = 7'h1F;

parameter ADDR_20 = 7'h20;
parameter ADDR_21 = 7'h21;
parameter ADDR_22 = 7'h22;
parameter ADDR_23 = 7'h23;
parameter ADDR_24 = 7'h24;
parameter ADDR_25 = 7'h25;
parameter ADDR_26 = 7'h26;
parameter ADDR_27 = 7'h27;
parameter ADDR_28 = 7'h28;
parameter ADDR_29 = 7'h29;
parameter ADDR_2A = 7'h2A;
parameter ADDR_2B = 7'h2B;
parameter ADDR_2C = 7'h2C;
parameter ADDR_2D = 7'h2D;
parameter ADDR_2E = 7'h2E;
parameter ADDR_2F = 7'h2F;

parameter ADDR_30 = 7'h30;
parameter ADDR_31 = 7'h31;
parameter ADDR_32 = 7'h32;
parameter ADDR_33 = 7'h33;
parameter ADDR_34 = 7'h34;
parameter ADDR_35 = 7'h35;
parameter ADDR_36 = 7'h36;
parameter ADDR_37 = 7'h37;
parameter ADDR_38 = 7'h38;
parameter ADDR_39 = 7'h39;
parameter ADDR_3A = 7'h3A;
parameter ADDR_3B = 7'h3B;
parameter ADDR_3C = 7'h3C;
parameter ADDR_3D = 7'h3D;
parameter ADDR_3E = 7'h3E;
parameter ADDR_3F = 7'h3F;

parameter ADDR_40 = 7'h40;
parameter ADDR_41 = 7'h41;
parameter ADDR_42 = 7'h42;
parameter ADDR_43 = 7'h43;
parameter ADDR_44 = 7'h44;
parameter ADDR_45 = 7'h45;
parameter ADDR_46 = 7'h46;
parameter ADDR_47 = 7'h47;
parameter ADDR_48 = 7'h48;
parameter ADDR_49 = 7'h49;
parameter ADDR_4A = 7'h4A;
parameter ADDR_4B = 7'h4B;
parameter ADDR_4C = 7'h4C;
parameter ADDR_4D = 7'h4D;
parameter ADDR_4E = 7'h4E;
parameter ADDR_4F = 7'h4F;

parameter ADDR_50 = 7'h50;
parameter ADDR_51 = 7'h51;
parameter ADDR_52 = 7'h52;
parameter ADDR_53 = 7'h53;
parameter ADDR_54 = 7'h54;
parameter ADDR_55 = 7'h55;
parameter ADDR_56 = 7'h56;
parameter ADDR_57 = 7'h57;
parameter ADDR_58 = 7'h58;
parameter ADDR_59 = 7'h59;
parameter ADDR_5A = 7'h5A;
parameter ADDR_5B = 7'h5B;
parameter ADDR_5C = 7'h5C;
parameter ADDR_5D = 7'h5D;
parameter ADDR_5E = 7'h5E;
parameter ADDR_5F = 7'h5F;

parameter ADDR_60 = 7'h60;
parameter ADDR_61 = 7'h61;
parameter ADDR_62 = 7'h62;
parameter ADDR_63 = 7'h63;
parameter ADDR_64 = 7'h64;
parameter ADDR_65 = 7'h65;
parameter ADDR_66 = 7'h66;
parameter ADDR_67 = 7'h67;
parameter ADDR_68 = 7'h68;
parameter ADDR_69 = 7'h69;
parameter ADDR_6A = 7'h6A;
parameter ADDR_6B = 7'h6B;
parameter ADDR_6C = 7'h6C;
parameter ADDR_6D = 7'h6D;
parameter ADDR_6E = 7'h6E;
parameter ADDR_6F = 7'h6F;

parameter ADDR_70 = 7'h70;
parameter ADDR_71 = 7'h71;
parameter ADDR_72 = 7'h72;
parameter ADDR_73 = 7'h73;
parameter ADDR_74 = 7'h74;
parameter ADDR_75 = 7'h75;
parameter ADDR_76 = 7'h76;
parameter ADDR_77 = 7'h77;
parameter ADDR_78 = 7'h78;
parameter ADDR_79 = 7'h79;
parameter ADDR_7A = 7'h7A;
parameter ADDR_7B = 7'h7B;
parameter ADDR_7C = 7'h7C;
parameter ADDR_7D = 7'h7D;
parameter ADDR_7E = 7'h7E;
parameter ADDR_7F = 7'h7F;

always @(*) begin
	case (addr)
		ADDR_00: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001;
		ADDR_01: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010;
		ADDR_02: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100;
		ADDR_03: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000;
		ADDR_04: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000;
		ADDR_05: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000;
		ADDR_06: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000;
		ADDR_07: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000;
		ADDR_08: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000;
		ADDR_09: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000;
		ADDR_0A: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000;
		ADDR_0B: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000;
		ADDR_0C: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000;
		ADDR_0D: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000;
		ADDR_0E: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000;
		ADDR_0F: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000;

		ADDR_10: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000;
		ADDR_11: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000;
		ADDR_12: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000;
		ADDR_13: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000;
		ADDR_14: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000;
		ADDR_15: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000;
		ADDR_16: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000;
		ADDR_17: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000;
		ADDR_18: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000;
		ADDR_19: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000;
		ADDR_1A: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000;
		ADDR_1B: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000;
		ADDR_1C: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000;
		ADDR_1D: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000;
		ADDR_1E: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000;
		ADDR_1F: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000;

		ADDR_20: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_21: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_22: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_23: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_24: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_25: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_26: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_27: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_28: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_29: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_2A: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_2B: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_2C: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_2D: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_2E: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_2F: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

		ADDR_30: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_31: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_32: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_33: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_34: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_35: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_36: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_37: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_38: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_39: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_3A: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_3B: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_3C: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_3D: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_3E: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_3F: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

		ADDR_40: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_41: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_42: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_43: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_44: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_45: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_46: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_47: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_48: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_49: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_4A: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_4B: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_4C: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_4D: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_4E: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_4F: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

		ADDR_50: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_51: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_52: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_53: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_54: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_55: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_56: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_57: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_58: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_59: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_5A: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_5B: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_5C: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_5D: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_5E: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_5F: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

		ADDR_60: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_61: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_62: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_63: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_64: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_65: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_66: reg_sel = 128'b0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_67: reg_sel = 128'b0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_68: reg_sel = 128'b0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_69: reg_sel = 128'b0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_6A: reg_sel = 128'b0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_6B: reg_sel = 128'b0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_6C: reg_sel = 128'b0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_6D: reg_sel = 128'b0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_6E: reg_sel = 128'b0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_6F: reg_sel = 128'b0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

		ADDR_70: reg_sel = 128'b0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_71: reg_sel = 128'b0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_72: reg_sel = 128'b0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_73: reg_sel = 128'b0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_74: reg_sel = 128'b0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_75: reg_sel = 128'b0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_76: reg_sel = 128'b0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_77: reg_sel = 128'b0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_78: reg_sel = 128'b0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_79: reg_sel = 128'b0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_7A: reg_sel = 128'b0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_7B: reg_sel = 128'b0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_7C: reg_sel = 128'b0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_7D: reg_sel = 128'b0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_7E: reg_sel = 128'b0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		ADDR_7F: reg_sel = 128'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
	endcase
end

assign wr_sel[0] = reg_sel[0] & wr_en;
assign wr_sel[1] = reg_sel[1] & wr_en;
assign wr_sel[2] = reg_sel[2] & wr_en;
assign wr_sel[3] = reg_sel[3] & wr_en;
assign wr_sel[4] = reg_sel[4] & wr_en;
assign wr_sel[5] = reg_sel[5] & wr_en;
assign wr_sel[6] = reg_sel[6] & wr_en;
assign wr_sel[7] = reg_sel[7] & wr_en;
assign wr_sel[8] = reg_sel[8] & wr_en;
assign wr_sel[9] = reg_sel[9] & wr_en;

assign wr_sel[10] = reg_sel[10] & wr_en;
assign wr_sel[11] = reg_sel[11] & wr_en;
assign wr_sel[12] = reg_sel[12] & wr_en;
assign wr_sel[13] = reg_sel[13] & wr_en;
assign wr_sel[14] = reg_sel[14] & wr_en;
assign wr_sel[15] = reg_sel[15] & wr_en;
assign wr_sel[16] = reg_sel[16] & wr_en;
assign wr_sel[17] = reg_sel[17] & wr_en;
assign wr_sel[18] = reg_sel[18] & wr_en;
assign wr_sel[19] = reg_sel[19] & wr_en;

assign wr_sel[20] = reg_sel[20] & wr_en;
assign wr_sel[21] = reg_sel[21] & wr_en;
assign wr_sel[22] = reg_sel[22] & wr_en;
assign wr_sel[23] = reg_sel[23] & wr_en;
assign wr_sel[24] = reg_sel[24] & wr_en;
assign wr_sel[25] = reg_sel[25] & wr_en;
assign wr_sel[26] = reg_sel[26] & wr_en;
assign wr_sel[27] = reg_sel[27] & wr_en;
assign wr_sel[28] = reg_sel[28] & wr_en;
assign wr_sel[29] = reg_sel[29] & wr_en;

assign wr_sel[30] = reg_sel[30] & wr_en;
assign wr_sel[31] = reg_sel[31] & wr_en;
assign wr_sel[32] = reg_sel[32] & wr_en;
assign wr_sel[33] = reg_sel[33] & wr_en;
assign wr_sel[34] = reg_sel[34] & wr_en;
assign wr_sel[35] = reg_sel[35] & wr_en;
assign wr_sel[36] = reg_sel[36] & wr_en;
assign wr_sel[37] = reg_sel[37] & wr_en;
assign wr_sel[38] = reg_sel[38] & wr_en;
assign wr_sel[39] = reg_sel[39] & wr_en;

assign wr_sel[40] = reg_sel[40] & wr_en;
assign wr_sel[41] = reg_sel[41] & wr_en;
assign wr_sel[42] = reg_sel[42] & wr_en;
assign wr_sel[43] = reg_sel[43] & wr_en;
assign wr_sel[44] = reg_sel[44] & wr_en;
assign wr_sel[45] = reg_sel[45] & wr_en;
assign wr_sel[46] = reg_sel[46] & wr_en;
assign wr_sel[47] = reg_sel[47] & wr_en;
assign wr_sel[48] = reg_sel[48] & wr_en;
assign wr_sel[49] = reg_sel[49] & wr_en;

assign wr_sel[50] = reg_sel[50] & wr_en;
assign wr_sel[51] = reg_sel[51] & wr_en;
assign wr_sel[52] = reg_sel[52] & wr_en;
assign wr_sel[53] = reg_sel[53] & wr_en;
assign wr_sel[54] = reg_sel[54] & wr_en;
assign wr_sel[55] = reg_sel[55] & wr_en;
assign wr_sel[56] = reg_sel[56] & wr_en;
assign wr_sel[57] = reg_sel[57] & wr_en;
assign wr_sel[58] = reg_sel[58] & wr_en;
assign wr_sel[59] = reg_sel[59] & wr_en;

assign wr_sel[60] = reg_sel[60] & wr_en;
assign wr_sel[61] = reg_sel[61] & wr_en;
assign wr_sel[62] = reg_sel[62] & wr_en;
assign wr_sel[63] = reg_sel[63] & wr_en;
assign wr_sel[64] = reg_sel[64] & wr_en;
assign wr_sel[65] = reg_sel[65] & wr_en;
assign wr_sel[66] = reg_sel[66] & wr_en;
assign wr_sel[67] = reg_sel[67] & wr_en;
assign wr_sel[68] = reg_sel[68] & wr_en;
assign wr_sel[69] = reg_sel[69] & wr_en;

assign wr_sel[70] = reg_sel[70] & wr_en;
assign wr_sel[71] = reg_sel[71] & wr_en;
assign wr_sel[72] = reg_sel[72] & wr_en;
assign wr_sel[73] = reg_sel[73] & wr_en;
assign wr_sel[74] = reg_sel[74] & wr_en;
assign wr_sel[75] = reg_sel[75] & wr_en;
assign wr_sel[76] = reg_sel[76] & wr_en;
assign wr_sel[77] = reg_sel[77] & wr_en;
assign wr_sel[78] = reg_sel[78] & wr_en;
assign wr_sel[79] = reg_sel[79] & wr_en;

assign wr_sel[80] = reg_sel[80] & wr_en;
assign wr_sel[81] = reg_sel[81] & wr_en;
assign wr_sel[82] = reg_sel[82] & wr_en;
assign wr_sel[83] = reg_sel[83] & wr_en;
assign wr_sel[84] = reg_sel[84] & wr_en;
assign wr_sel[85] = reg_sel[85] & wr_en;
assign wr_sel[86] = reg_sel[86] & wr_en;
assign wr_sel[87] = reg_sel[87] & wr_en;
assign wr_sel[88] = reg_sel[88] & wr_en;
assign wr_sel[89] = reg_sel[89] & wr_en;

assign wr_sel[90] = reg_sel[90] & wr_en;
assign wr_sel[91] = reg_sel[91] & wr_en;
assign wr_sel[92] = reg_sel[92] & wr_en;
assign wr_sel[93] = reg_sel[93] & wr_en;
assign wr_sel[94] = reg_sel[94] & wr_en;
assign wr_sel[95] = reg_sel[95] & wr_en;
assign wr_sel[96] = reg_sel[96] & wr_en;
assign wr_sel[97] = reg_sel[97] & wr_en;
assign wr_sel[98] = reg_sel[98] & wr_en;
assign wr_sel[99] = reg_sel[99] & wr_en;

assign wr_sel[100] = reg_sel[100] & wr_en;
assign wr_sel[101] = reg_sel[101] & wr_en;
assign wr_sel[102] = reg_sel[102] & wr_en;
assign wr_sel[103] = reg_sel[103] & wr_en;
assign wr_sel[104] = reg_sel[104] & wr_en;
assign wr_sel[105] = reg_sel[105] & wr_en;
assign wr_sel[106] = reg_sel[106] & wr_en;
assign wr_sel[107] = reg_sel[107] & wr_en;
assign wr_sel[108] = reg_sel[108] & wr_en;
assign wr_sel[109] = reg_sel[109] & wr_en;

assign wr_sel[110] = reg_sel[110] & wr_en;
assign wr_sel[111] = reg_sel[111] & wr_en;
assign wr_sel[112] = reg_sel[112] & wr_en;
assign wr_sel[113] = reg_sel[113] & wr_en;
assign wr_sel[114] = reg_sel[114] & wr_en;
assign wr_sel[115] = reg_sel[115] & wr_en;
assign wr_sel[116] = reg_sel[116] & wr_en;
assign wr_sel[117] = reg_sel[117] & wr_en;
assign wr_sel[118] = reg_sel[118] & wr_en;
assign wr_sel[119] = reg_sel[119] & wr_en;

assign wr_sel[120] = reg_sel[120] & wr_en;
assign wr_sel[121] = reg_sel[121] & wr_en;
assign wr_sel[122] = reg_sel[122] & wr_en;
assign wr_sel[123] = reg_sel[123] & wr_en;
assign wr_sel[124] = reg_sel[124] & wr_en;
assign wr_sel[125] = reg_sel[125] & wr_en;
assign wr_sel[126] = reg_sel[126] & wr_en;
assign wr_sel[127] = reg_sel[127] & wr_en;

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_00 <= 9'b001001000;
	else if (wr_sel[0] == 1)
		addr_00 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_01 <= 9'b000000001;
	else if (wr_sel[1] == 1)
		addr_01 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_02 <= 9'b001010000;
	else if (wr_sel[2] == 1)
		addr_02 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_03 <= 9'b000000000;
	else if (wr_sel[3] == 1)
		addr_03 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_04 <= 9'b001011000;
	else if (wr_sel[4] == 1)
		addr_04 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_05 <= 9'b010000000;
	else if (wr_sel[5] == 1)
		addr_05 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_06 <= 9'b101010011;
	else if (wr_sel[6] == 1)
		addr_06 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_07 <= 9'b010010001;
	else if (wr_sel[7] == 1)
		addr_07 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_08 <= 9'b001011000;
	else if (wr_sel[8] == 1)
		addr_08 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_09 <= 9'b111111111;
	else if (wr_sel[9] == 1)
		addr_09 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_0a <= 9'b000101111;
	else if (wr_sel[10] == 1)
		addr_0a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_0b <= 9'b001100000;
	else if (wr_sel[11] == 1)
		addr_0b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_0c <= 9'b111111111;
	else if (wr_sel[12] == 1)
		addr_0c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_0d <= 9'b000000111;
	else if (wr_sel[13] == 1)
		addr_0d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_0e <= 9'b011100001;
	else if (wr_sel[14] == 1)
		addr_0e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_0f <= 9'b110111000;
	else if (wr_sel[15] == 1)
		addr_0f <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_10 <= 9'b011011001;
	else if (wr_sel[16] == 1)
		addr_10 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_11 <= 9'b110111101;
	else if (wr_sel[17] == 1)
		addr_11 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_12 <= 9'b001111000;
	else if (wr_sel[18] == 1)
		addr_12 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n)
		addr_13 <= 9'b000000100;
	else if (wr_sel[19] == 1)
		addr_13 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n) 
		addr_14 <= 9'b000000000;
	else if (wr_sel[20] == 1) 
		addr_14 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin
	if (!rst_n) 
		addr_15 <= 9'b000000000;
	else if (wr_sel[21] == 1) 
		addr_15 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_16 <= 9'b000000000;
	else if (wr_sel[22] == 1) 
		addr_16 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_17 <= 9'b000000000;
	else if (wr_sel[23] == 1) 
		addr_17 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_18 <= 9'b000000000;
	else if (wr_sel[24] == 1) 
		addr_18 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_19 <= 9'b000000000;
	else if (wr_sel[25] == 1) 
		addr_19 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_1a <= 9'b000000000;
	else if (wr_sel[26] == 1) 
		addr_1a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_1b <= 9'b000000000;
	else if (wr_sel[27] == 1) 
		addr_1b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_1c <= 9'b000000000;
	else if (wr_sel[28] == 1) 
		addr_1c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_1d <= 9'b000000000;
	else if (wr_sel[29] == 1) 
		addr_1d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_1e <= 9'b000000000;
	else if (wr_sel[30] == 1) 
		addr_1e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_1f <= 9'b000000000;
	else if (wr_sel[31] == 1) 
		addr_1f <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_20 <= 9'b000000000;
	else if (wr_sel[32] == 1) 
		addr_20 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_21 <= 9'b000000000;
	else if (wr_sel[33] == 1) 
		addr_21 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_22 <= 9'b000000000;
	else if (wr_sel[34] == 1) 
		addr_22 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_23 <= 9'b000000000;
	else if (wr_sel[35] == 1) 
		addr_23 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_24 <= 9'b000000000;
	else if (wr_sel[36] == 1) 
		addr_24 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_25 <= 9'b000000000;
	else if (wr_sel[37] == 1) 
		addr_25 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_26 <= 9'b000000000;
	else if (wr_sel[38] == 1) 
		addr_26 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_27 <= 9'b000000000;
	else if (wr_sel[39] == 1) 
		addr_27 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_28 <= 9'b000000000;
	else if (wr_sel[40] == 1) 
		addr_28 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_29 <= 9'b000000000;
	else if (wr_sel[41] == 1) 
		addr_29 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_2a <= 9'b000000000;
	else if (wr_sel[42] == 1) 
		addr_2a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_2b <= 9'b000000000;
	else if (wr_sel[43] == 1) 
		addr_2b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_2c <= 9'b000000000;
	else if (wr_sel[44] == 1) 
		addr_2c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_2d <= 9'b000000000;
	else if (wr_sel[45] == 1) 
		addr_2d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_2e <= 9'b000000000;
	else if (wr_sel[46] == 1) 
		addr_2e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_2f <= 9'b000000000;
	else if (wr_sel[47] == 1) 
		addr_2f <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_30 <= 9'b000000000;
	else if (wr_sel[48] == 1) 
		addr_30 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_31 <= 9'b000000000;
	else if (wr_sel[49] == 1) 
		addr_31 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_32 <= 9'b000000000;
	else if (wr_sel[50] == 1) 
		addr_32 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_33 <= 9'b000000000;
	else if (wr_sel[51] == 1) 
		addr_33 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_34 <= 9'b000000000;
	else if (wr_sel[52] == 1) 
		addr_34 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_35 <= 9'b000000000;
	else if (wr_sel[53] == 1) 
		addr_35 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_36 <= 9'b000000000;
	else if (wr_sel[54] == 1) 
		addr_36 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_37 <= 9'b000000000;
	else if (wr_sel[55] == 1) 
		addr_37 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_38 <= 9'b000000000;
	else if (wr_sel[56] == 1) 
		addr_38 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_39 <= 9'b000000000;
	else if (wr_sel[57] == 1) 
		addr_39 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_3a <= 9'b000000000;
	else if (wr_sel[58] == 1) 
		addr_3a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_3b <= 9'b000000000;
	else if (wr_sel[59] == 1) 
		addr_3b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_3c <= 9'b000000000;
	else if (wr_sel[60] == 1) 
		addr_3c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_3d <= 9'b000000000;
	else if (wr_sel[61] == 1) 
		addr_3d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_3e <= 9'b000000000;
	else if (wr_sel[62] == 1) 
		addr_3e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_3f <= 9'b000000000;
	else if (wr_sel[63] == 1) 
		addr_3f <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_40 <= 9'b000000000;
	else if (wr_sel[64] == 1) 
		addr_40 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_41 <= 9'b000000000;
	else if (wr_sel[65] == 1) 
		addr_41 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_42 <= 9'b000000000;
	else if (wr_sel[66] == 1) 
		addr_42 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_43 <= 9'b000000000;
	else if (wr_sel[67] == 1) 
		addr_43 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_44 <= 9'b000000000;
	else if (wr_sel[68] == 1) 
		addr_44 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_45 <= 9'b000000000;
	else if (wr_sel[69] == 1) 
		addr_45 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_46 <= 9'b000000000;
	else if (wr_sel[70] == 1) 
		addr_46 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_47 <= 9'b000000000;
	else if (wr_sel[71] == 1) 
		addr_47 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_48 <= 9'b000000000;
	else if (wr_sel[72] == 1) 
		addr_48 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_49 <= 9'b000000000;
	else if (wr_sel[73] == 1) 
		addr_49 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_4a <= 9'b000000000;
	else if (wr_sel[74] == 1) 
		addr_4a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_4b <= 9'b000000000;
	else if (wr_sel[75] == 1) 
		addr_4b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_4c <= 9'b000000000;
	else if (wr_sel[76] == 1) 
		addr_4c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_4d <= 9'b000000000;
	else if (wr_sel[77] == 1) 
		addr_4d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_4e <= 9'b000000000;
	else if (wr_sel[78] == 1) 
		addr_4e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_4f <= 9'b000000000;
	else if (wr_sel[79] == 1) 
		addr_4f <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_50 <= 9'b000000000;
	else if (wr_sel[80] == 1) 
		addr_50 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_51 <= 9'b000000000;
	else if (wr_sel[81] == 1) 
		addr_51 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_52 <= 9'b000000000;
	else if (wr_sel[82] == 1) 
		addr_52 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_53 <= 9'b000000000;
	else if (wr_sel[83] == 1) 
		addr_53 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_54 <= 9'b000000000;
	else if (wr_sel[84] == 1) 
		addr_54 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_55 <= 9'b000000000;
	else if (wr_sel[85] == 1) 
		addr_55 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_56 <= 9'b000000000;
	else if (wr_sel[86] == 1) 
		addr_56 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_57 <= 9'b000000000;
	else if (wr_sel[87] == 1) 
		addr_57 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_58 <= 9'b000000000;
	else if (wr_sel[88] == 1) 
		addr_58 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_59 <= 9'b000000000;
	else if (wr_sel[89] == 1) 
		addr_59 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_5a <= 9'b000000000;
	else if (wr_sel[90] == 1) 
		addr_5a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_5b <= 9'b000000000;
	else if (wr_sel[91] == 1) 
		addr_5b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_5c <= 9'b000000000;
	else if (wr_sel[92] == 1) 
		addr_5c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_5d <= 9'b000000000;
	else if (wr_sel[93] == 1) 
		addr_5d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_5e <= 9'b000000000;
	else if (wr_sel[94] == 1) 
		addr_5e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_5f <= 9'b000000000;
	else if (wr_sel[95] == 1) 
		addr_5f <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_60 <= 9'b000000000;
	else if (wr_sel[96] == 1) 
		addr_60 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_61 <= 9'b000000000;
	else if (wr_sel[97] == 1) 
		addr_61 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_62 <= 9'b000000000;
	else if (wr_sel[98] == 1) 
		addr_62 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_63 <= 9'b000000000;
	else if (wr_sel[99] == 1) 
		addr_63 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_64 <= 9'b000000000;
	else if (wr_sel[100] == 1) 
		addr_64 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_65 <= 9'b000000000;
	else if (wr_sel[101] == 1) 
		addr_65 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_66 <= 9'b000000000;
	else if (wr_sel[102] == 1) 
		addr_66 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_67 <= 9'b000000000;
	else if (wr_sel[103] == 1) 
		addr_67 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_68 <= 9'b000000000;
	else if (wr_sel[104] == 1) 
		addr_68 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_69 <= 9'b000000000;
	else if (wr_sel[105] == 1) 
		addr_69 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_6a <= 9'b000000000;
	else if (wr_sel[106] == 1) 
		addr_6a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_6b <= 9'b000000000;
	else if (wr_sel[107] == 1) 
		addr_6b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_6c <= 9'b000000000;
	else if (wr_sel[108] == 1) 
		addr_6c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_6d <= 9'b000000000;
	else if (wr_sel[109] == 1) 
		addr_6d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_6e <= 9'b000000000;
	else if (wr_sel[110] == 1) 
		addr_6e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_6f <= 9'b000000000;
	else if (wr_sel[111] == 1) 
		addr_6f <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_70 <= 9'b000000000;
	else if (wr_sel[112] == 1) 
		addr_70 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_71 <= 9'b000000000;
	else if (wr_sel[113] == 1) 
		addr_71 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_72 <= 9'b000000000;
	else if (wr_sel[114] == 1) 
		addr_72 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_73 <= 9'b000000000;
	else if (wr_sel[115] == 1) 
		addr_73 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_74 <= 9'b000000000;
	else if (wr_sel[116] == 1) 
		addr_74 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_75 <= 9'b000000000;
	else if (wr_sel[117] == 1) 
		addr_75 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_76 <= 9'b000000000;
	else if (wr_sel[118] == 1) 
		addr_76 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_77 <= 9'b000000000;
	else if (wr_sel[119] == 1) 
		addr_77 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_78 <= 9'b000000000;
	else if (wr_sel[120] == 1) 
		addr_78 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_79 <= 9'b000000000;
	else if (wr_sel[121] == 1) 
		addr_79 <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_7a <= 9'b000000000;
	else if (wr_sel[122] == 1) 
		addr_7a <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_7b <= 9'b000000000;
	else if (wr_sel[123] == 1) 
		addr_7b <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_7c <= 9'b000000000;
	else if (wr_sel[124] == 1) 
		addr_7c <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_7d <= 9'b000000000;
	else if (wr_sel[125] == 1) 
		addr_7d <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_7e <= 9'b000000000;
	else if (wr_sel[126] == 1) 
		addr_7e <= data[8:0];
end

always @(posedge clk or negedge rst_n) begin 
	if (!rst_n) 
		addr_7f <= 9'b000000000;
	else if (wr_sel[127] == 1) 
		addr_7f <= data[8:0];
end

always @(*) begin
	case (reg_sel)

		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001: q = addr_00;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010: q = addr_01;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100: q = addr_02;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000: q = addr_03;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000: q = addr_04;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000: q = addr_05;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000: q = addr_06;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000: q = addr_07;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000: q = addr_08;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000: q = addr_09;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000: q = addr_0a;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000: q = addr_0b;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000: q = addr_0c;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000: q = addr_0d;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000: q = addr_0e;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000: q = addr_0f;

		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000: q = addr_10;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000: q = addr_11;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000: q = addr_12;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000: q = addr_13;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000: q = addr_14;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000: q = addr_15;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000: q = addr_16;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000: q = addr_17;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000: q = addr_18;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000: q = addr_19;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000: q = addr_1a;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000: q = addr_1b;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000: q = addr_1c;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000: q = addr_1d;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000: q = addr_1e;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000: q = addr_1f;

		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_20;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_21;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_22;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_23;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_24;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_25;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_26;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_27;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_28;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_29;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_2a;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_2b;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_2c;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_2d;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_2e;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_2f;

		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_30;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_31;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_32;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_33;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_34;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_35;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_36;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_37;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_38;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_39;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_3a;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_3b;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_3c;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_3d;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_3e;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_3f;

		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_40;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_41;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_42;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_43;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_44;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_45;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_46;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_47;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_48;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_49;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_4a;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_4b;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_4c;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_4d;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_4e;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_4f;

		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_50;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_51;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_52;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_53;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_54;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_55;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_56;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_57;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_58;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_59;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_5a;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_5b;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_5c;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_5d;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_5e;
		128'b0000_0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_5f;

		128'b0000_0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_60;
		128'b0000_0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_61;
		128'b0000_0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_62;
		128'b0000_0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_63;
		128'b0000_0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_64;
		128'b0000_0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_65;
		128'b0000_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_66;
		128'b0000_0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_67;
		128'b0000_0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_68;
		128'b0000_0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_69;
		128'b0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_6a;
		128'b0000_0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_6b;
		128'b0000_0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_6c;
		128'b0000_0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_6d;
		128'b0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_6e;
		128'b0000_0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_6f;

		128'b0000_0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_70;
		128'b0000_0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_71;
		128'b0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_72;
		128'b0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_73;
		128'b0000_0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_74;
		128'b0000_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_75;
		128'b0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_76;
		128'b0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_77;
		128'b0000_0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_78;
		128'b0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_79;
		128'b0000_0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_7a;
		128'b0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_7b;
		128'b0001_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_7c;
		128'b0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_7d;
		128'b0100_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_7e;
		128'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000: q = addr_7f;

		default: q = 9'b0;

	endcase
end
endmodule
